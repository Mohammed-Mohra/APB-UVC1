`include "example_test.svh"
