`include "moh_apb_if.sv"

package moh_apb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  typedef uvm_config_db#(virtual moh_apb_if) apb_vif_config;

  `include "moh_apb_types.svh"
  `include "moh_apb_config_class.sv"
  `include "moh_apb_seq_item.sv"

  // Requester files
  `include "moh_apb_requester_sequence_lib.sv"
  `include "moh_apb_monitor.sv"
  `include "moh_apb_requester_sequencer.sv"
  `include "moh_apb_requester_driver.sv"
  `include "moh_apb_requester_agent.sv"

  //Completer files
  `include "moh_apb_completer_sequencer.sv"
  `include "moh_apb_completer_sequence_lib.sv"
  `include "moh_apb_completer_driver.sv"
  `include "moh_apb_completer_agent.sv"
  `include "moh_apb_env.sv"

endpackage : moh_apb_pkg
