`ifndef __MOH_APB_EXAMPLE_PKG_SV
`define __MOH_APB_EXAMPLE_PKG_SV

package moh_apb_example_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  import moh_apb_pkg::*;

  `include "moh_apb_virtual_sequencer.sv"
  `include "moh_apb_virtual_sequence.sv"
  `include "moh_apb_example_env.sv"
  `include "moh_apb_base_test.sv"
  `include "uvm_test_lib.sv"
endpackage : moh_apb_example_pkg

`endif
